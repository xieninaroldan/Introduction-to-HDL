module Group3_Lab4_full(A,B,Bin,Diff,Bout);
input A,B,Bin;
output Diff,Bout;

endmodule