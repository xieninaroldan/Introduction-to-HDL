module Group3_Lab3(a1,a2,a3,b);
input a1,a2,a3;
output b;

endmodule