module Group3_Lab4(a1,a2,b,b1,b2);
input a1,a2,b2;
output b,b1;

endmodule